.OPTION LIMPTS = 501


VDD 4 0 DC 2.5 AC 1.0
VSS 0 5 DC 2.5


* solve   2x + 3y = 40
*         2x + y  = 5

* begin
xamp1 inp inm out 4 5  opamp
rf inm out 100k
r1 out2 inm 66.7k


rpf inp  0 100k

Vcoeff  vrp1 0 dc 2

*VDCfromop vfrom 0 dc 2
*xtest vrp1 out settling_test v0=0 v1=2 interval=10u

rp1  vrp1 inp 100k

rpy  inp 0 200k
* end

* opamp for Y coordinate
* begin
xamp2 inp2 inm2 out2 4 5  opamp
rf2 inm2 out2 100k
r12 out inm2 50k


rpf2 inp2  0 100k

Vcoeff2  vrp2 0 dc 0.5 

*xtest2 vrp2 out2 settling_test v0=0 v1=0.5 interval=10u

rp12  vrp2 inp2 100k

rpy2  inp2 0 100k

.subckt opamp 1 2 6 8 9

M1 4 2 3 3 NMOS1 W = 3U L = 1U AD = 18P AS = 18P PD = 18U PS = 18U
M2 5 1 3 3 NMOS1 W = 3U L = 1U AD = 18P AS = 18P PD = 18U PS = 18U
M3 4 4 8 8 PMOS1 W = 15U L = 1U AD = 90P AS = 90P PD = 42U PS = 42U
M4 5 4 8 8 PMOS1 W = 15U L = 1U AD = 90P AS = 90P PD = 42U PS = 42U

M5 3 7 9 9 NMOS1 W = 4.5U L = 1U AD = 27P AS = 27P PD = 21U PS = 21U

M6 6 5 8 8 PMOS1 W = 94U L = 1U AD = 564P AS = 564P PD = 200U PS = 200U

M7 6 7 9 9 NMOS1 W = 14U L = 1U AD = 84P AS = 84P PD = 40U PS = 40U

M8 7 7 9 9 NMOS1 W = 4.5U L = 1U AD = 27P AS = 27P PD = 21U PS = 21U

CC 5 6 3.0P

.MODEL NMOS1 NMOS VTO = 0.70 KP = 110U GAMMA = 0.4  LAMBDA = 0.04 PHI =
+ 0.7 MJ = 0.5 MJSW = 0.38  CGBO = 700P  CGSO = 220P CGDO = 220P CJ
+ = 770U CJSW = 380P LD = 0.016U TOX = 14N

.MODEL PMOS1 PMOS VTO = -0.70 KP = 50U GAMMA = 0.57  LAMBDA = 0.05 PHI =
+ 0.8 MJ = 0.5 MJSW = 0.35  CGBO = 700P  CGSO = 220P CGDO = 220P CJ
+ = 560U CJSW = 350P LD = 0.014U TOX = 14N

IBIAS 8 7 30U

.ENDS


* end

*.DC Vcoeff -1 20 0.1
*.DC Vcoeff2 -1 5 0.1

* Correct out = -0.625V   out2=1.75V
.PROBE V(out)
.PROBE V(out2)

* diverges if simulated for more than 4u
.tran 10p 6u 0.0 0.01u

***--------------------------
.OPTION  INGOLD=2 ARTIST=2 PSF=2 PROBE=0 GMMIN=1e-15 METHOD=GEAR
.OPTION POST
*.TEMP  30
.OPTIONS SCALE = 1.00
.SAVE

.end
